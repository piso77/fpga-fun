// CPU opcodes

`define ADD_OP 4'b0000
`define SUB_OP 4'b0001
`define MUL_OP 4'b0010
`define SHL_OP 4'b0011
`define SHR_OP 4'b0100
`define ROL_OP 4'b0101
`define ROR_OP 4'b0110
`define OR_OP  4'b0111
`define AND_OP 4'b1000
`define XOR_OP 4'b1001
`define LDI_OP 4'b1010
`define LDR_OP 4'b1011
`define MV_OP  4'b1100
`define ST_OP  4'b1101
`define BRI_OP 4'b1110
`define BRR_OP 4'b1111
