/*
Displays a grid of digits on the CRT using a RAM module.
*/

module ram_text_top(clk, reset, hsync, vsync, rgb);
input clk, reset;
output hsync, vsync;
output [2:0] rgb;



endmodule
